module displayEncoder(
	// TODO: define your input and output ports
	
);
	// TODO: create signals for the six 4-bit digits
	
	// TODO: Instantiate six copies of sevenSegDigit, one for each digit (calculated below) 

	// The following block contains the logic of your combinational circuit
	always_comb begin
		// TODO: Convert a 20-bit input result to six individual digits (4 bits each) 

	end

endmodule