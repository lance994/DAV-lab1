//module sevenSegDigit(
	// TODO: define your input and output ports

//);

	// The following block contains the logic of your combinational circuit
	//always_comb begin
		// TODO: fill out the case construct below to output the correct seven-segment display bits
		//case (/* */)
			
			//default: begin // this is the "catch-all" case - if none of the above cases match, this will execute
				/* TODO: set your output bits */

			//end
//		endcase
	//end

//endmodule
